//First module

module my_module(
    input logic a, b,
    output logic o
);
    assign o = a & b;

endmodule