//First module

module my_module(
    input logic a, b,
    output logic o
)
    and(o, a, b);

endmodule